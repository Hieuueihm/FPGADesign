LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_unsigned.ALL;

ENTITY Read_Pointer IS
    GENERIC (
        ADDR_WIDTH : INTEGER := 4
    );
    PORT (
        clk : IN STD_LOGIC;
        rd : IN STD_LOGIC;
        base_addr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
        fifo_empty : IN STD_LOGIC;
        fifo_re : OUT STD_LOGIC;
        rptr : OUT STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0)
    );
END ENTITY Read_Pointer;
ARCHITECTURE behavioral OF Read_Pointer IS
    SIGNAL read_addr : STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
    SIGNAL re : STD_LOGIC;
    SIGNAL initialized : BOOLEAN := FALSE; -- To track initialization state

BEGIN
    re <= (NOT fifo_empty) AND rd;
    fifo_re <= re;
    rptr <= read_addr;
    PROCESS (clk)
    BEGIN
        IF (rising_edge(clk)) THEN
            IF (NOT initialized) THEN
                read_addr <= base_addr;
                initialized <= TRUE;
            ELSIF (re = '1') THEN
                read_addr <= read_addr + STD_LOGIC_VECTOR(UNSIGNED(TO_UNSIGNED(1, ADDR_WIDTH)));
            END IF;
        END IF;
    END PROCESS;
END ARCHITECTURE behavioral;