`timescale 1ns / 1ps
module mips_top_tb (
    ports
);

endmodule
