LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
ENTITY DFF IS
    PORT (
        CLK : IN STD_LOGIC;
        EN : IN STD_LOGIC;
        D : IN STD_LOGIC;
        Q : OUT STD_LOGIC
    );
END ENTITY DFF;

ARCHITECTURE rtl OF DFF IS

BEGIN
    PROCESS (CLK)
    BEGIN
        IF rising_edge(CLK) THEN
            IF (en = '1') THEN
                Q <= D;
            END IF;
        END IF;
    END PROCESS;
END ARCHITECTURE rtl;