module moduleName (
    input clk,
    input [5:0] A1,A2, A3; // address of source and destination
    

);
    
endmodule