LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE STD.textio.ALL;

ENTITY ReadImage IS

    GENERIC (
        ADDR_WIDTH : INTEGER := 4;
        DATA_WIDTH : INTEGER := 8;
        IMAGE_SIZE : INTEGER := 15;
        IMAGE_FILE_NAME : STRING := "IMAGE_FILE.MIF"
    );
    PORT (
        clk : IN STD_LOGIC;
        data : IN STD_LOGIC_VECTOR((DATA_WIDTH - 1) DOWNTO 0);
        read_addr : IN STD_LOGIC_VECTOR((ADDR_WIDTH - 1) DOWNTO 0);
        write_addr : IN STD_LOGIC_VECTOR((ADDR_WIDTH - 1) DOWNTO 0);
        write_en : IN STD_LOGIC;
        read_en : IN STD_LOGIC;
        Q : OUT STD_LOGIC_VECTOR((DATA_WIDTH - 1) DOWNTO 0)
    );
END ENTITY ReadImage;
ARCHITECTURE behavioral OF ReadImage IS
    TYPE mem_type IS ARRAY(0 TO IMAGE_SIZE) OF STD_LOGIC_VECTOR((DATA_WIDTH - 1) DOWNTO 0);

    IMPURE FUNCTION init_mem(mif_file_name : IN STRING) RETURN mem_type IS
        FILE mif_file : text OPEN read_mode IS mif_file_name;
        VARIABLE mif_line : line;
        VARIABLE temp_bv : bit_vector(DATA_WIDTH - 1 DOWNTO 0);
        VARIABLE temp_mem : mem_type;

    BEGIN
        FOR i IN mem_type'RANGE LOOP
            readline(mif_file, mif_line);
            read(mif_line, temp_bv);
            temp_mem(i) := to_stdlogicvector(temp_bv);
        END LOOP;
        RETURN temp_mem;
    END FUNCTION;

    SIGNAL ram_block : mem_type := init_mem(IMAGE_FILE_NAME);
    SIGNAL read_address_reg : STD_LOGIC_VECTOR((ADDR_WIDTH - 1) DOWNTO 0) := (OTHERS => '0');

BEGIN
    PROCESS (clk)
    BEGIN
        IF (rising_edge(clk)) THEN
            IF (write_en = '1') THEN
                ram_block(to_integer(unsigned(write_addr))) <= data;
            END IF;
            IF (read_en = '1') THEN
                Q <= ram_block(to_integer(unsigned(read_addr)));
            END IF;
        END IF;
    END PROCESS;

END ARCHITECTURE behavioral;