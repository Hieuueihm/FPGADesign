LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
ENTITY UART_TX IS
    GENERIC (
        SYSTEM_CLK : INTEGER := 50_000_000;
        BAUD_RATE : INTEGER := 9_600;
        OS_RATE : INTEGER := 16;
        N : INTEGER := 8
    );
    PORT (
        CLK, RST : IN STD_LOGIC;
        Tx_start : IN STD_LOGIC;
        Tx_data_in : IN STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
        Tx_data_out : OUT STD_LOGIC;
        Tx_busy : OUT STD_LOGIC;
        Tx_finish : OUT STD_LOGIC
    );
END ENTITY UART_TX;

ARCHITECTURE rtl OF UART_TX IS
    CONSTANT CLK_BAUDRATE : INTEGER := SYSTEM_CLK / BAUD_RATE / OS_RATE;
    TYPE FSM IS(IDLE, START, DATA, STOP_S);
    SIGNAL STATE : FSM;
    SIGNAL tx_count : INTEGER RANGE 0 TO N - 1;
    SIGNAL count_clk : INTEGER RANGE 0 TO (CLK_BAUDRATE - 1);
    SIGNAL Tx_in : STD_LOGIC_VECTOR(N - 1 DOWNTO 0);
    SIGNAL Tx_out : STD_LOGIC;
    SIGNAL Tx_active : STD_LOGIC;
    SIGNAL Tx_end : STD_LOGIC;
BEGIN
    PROCESS (CLK, RST)

    BEGIN
        IF (RST = '1') THEN
            tx_count <= 0;
            count_clk <= 0;
            STATE <= IDLE;
            Tx_out <= '1';
            Tx_active <= '0';
            Tx_end <= '0';

        ELSIF (RISING_EDGE(CLK)) THEN
            CASE STATE IS
                WHEN IDLE =>
                    Tx_out <= '1';
                    Tx_active <= '0';
                    Tx_end <= '0';
                    count_clk <= 0;
                    tx_count <= 0;

                    IF (Tx_start = '1') THEN
                        Tx_in <= Tx_data_in;
                        STATE <= START;

                    ELSE
                        STATE <= IDLE;
                    END IF;
                WHEN START =>
                    Tx_out <= '0';
                    Tx_active <= '1'; --- activate Tx

                    IF (count_clk < (CLK_BAUDRATE - 1)) THEN
                        count_clk <= count_clk + 1;
                        STATE <= START;
                    ELSE
                        count_clk <= 0;
                        STATE <= DATA;
                    END IF;
                WHEN DATA =>
                    Tx_out <= Tx_in(tx_count);
                    IF (count_clk < (CLK_BAUDRATE - 1)) THEN
                        count_clk <= count_clk + 1;
                        STATE <= DATA;
                    ELSE
                        count_clk <= 0;
                        IF (tx_count < N - 1) THEN
                            tx_count <= tx_count + 1;
                            STATE <= DATA;
                        ELSE
                            tx_count <= 0;
                            STATE <= STOP_S;
                        END IF;
                    END IF;

                WHEN STOP_S =>

                    Tx_out <= '1';
                    IF (count_clk < (CLK_BAUDRATE - 1)) THEN
                        count_clk <= count_clk + 1;
                        STATE <= STOP_S;
                    ELSE
                        count_clk <= 0;
                        Tx_end <= '1';
                        Tx_active <= '0';
                        STATE <= IDLE;

                    END IF;

            END CASE;
        END IF;

    END PROCESS;
    Tx_data_out <= Tx_out;
    Tx_busy <= Tx_active;
    Tx_finish <= Tx_end;
END ARCHITECTURE rtl;