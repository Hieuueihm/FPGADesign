LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
ENTITY ALU IS

    PORT (
        A_BUS : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        B_BUS : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        ALU_ctrl : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- 4 bit
        ALU_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY ALU;
ARCHITECTURE rtl OF ALU IS

BEGIN

END ARCHITECTURE rtl;