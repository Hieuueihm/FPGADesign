LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
PACKAGE MyLib IS
    COMPONENT Read_Pointer IS
        GENERIC (
            ADDR_WIDTH : INTEGER := 4
        );
        PORT (
            clk : IN STD_LOGIC;
            rd : IN STD_LOGIC;
            -- fifo_empty : IN STD_LOGIC;
            base_addr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            fifo_re : OUT STD_LOGIC;

            rptr : OUT STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT Write_Pointer IS
        GENERIC (
            ADDR_WIDTH : INTEGER := 4
        );
        PORT (
            clk : IN STD_LOGIC;
            -- fifo_full : IN STD_LOGIC;
            wr : IN STD_LOGIC;
            base_addr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);

            wptr : OUT STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            fifo_we : OUT STD_LOGIC
        );
    END COMPONENT;
    COMPONENT Memory_Array IS
        GENERIC (
            ADDR_WIDTH : INTEGER := 4;
            DATA_WIDTH : INTEGER := 8
        );
        PORT (
            clk : IN STD_LOGIC;
            fifo_re : IN STD_LOGIC;
            fifo_we : IN STD_LOGIC;
            rptr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            wptr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            data_in : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
            data_out : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
        );
    END COMPONENT;
    COMPONENT Fifo_Memory IS

        GENERIC (
            ADDR_WIDTH : INTEGER := 4;
            DATA_WIDTH : INTEGER := 8
        );
        PORT (
            data_in : IN STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0);
            wr : IN STD_LOGIC;
            rd : IN STD_LOGIC;
            clk : IN STD_LOGIC;
            base_addr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            data_out : OUT STD_LOGIC_VECTOR(DATA_WIDTH - 1 DOWNTO 0)
        );
    END COMPONENT;

    COMPONENT Controller IS
        GENERIC (
            ADDR_WIDTH : INTEGER := 4
        );
        PORT (
            clk : IN STD_LOGIC;
            fifo_we : IN STD_LOGIC;
            fifo_rd : IN STD_LOGIC;
            wptr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            rptr : IN STD_LOGIC_VECTOR(ADDR_WIDTH - 1 DOWNTO 0);
            fifo_full : OUT STD_LOGIC;
            fifo_empty : OUT STD_LOGIC
        );
    END COMPONENT;
END PACKAGE MyLib;